------------------------------
-- Weicheng Huang            
-- testbench for lab
------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.components.all;

entity calculator_tb is
end calculator_tb;

architecture testbench of calculator_tb is
    -- Constants
    constant CLK_PERIOD : time := 20 ns; -- 50 MHz clock
    
    -- Signals
    signal clk          : std_logic := '0';
    signal reset        : std_logic := '1';
    signal reset_n      : std_logic := '0';
    signal execute      : std_logic := '0';
    signal ms           : std_logic := '0';
    signal mr           : std_logic := '0';
    signal switch       : std_logic_vector(7 downto 0) := (others => '0');
    signal op           : std_logic_vector(1 downto 0) := (others => '0');
    signal led          : std_logic_vector(3 downto 0);
    signal bcd_0        : std_logic_vector(6 downto 0);
    signal bcd_1        : std_logic_vector(6 downto 0);
    signal bcd_2        : std_logic_vector(6 downto 0);
    
    -- Test bench control
    signal test_complete : boolean := false;
    
    -- Component declaration
    component top
        port (
            clk       : in std_logic;
            reset_n   : in std_logic;
            execute   : in std_logic;
            ms        : in std_logic;
            mr        : in std_logic;
            switch    : in std_logic_vector(7 downto 0);
            op        : in std_logic_vector(1 downto 0);
            led       : out std_logic_vector(3 downto 0);
            bcd_0     : out std_logic_vector(6 downto 0);
            bcd_1     : out std_logic_vector(6 downto 0);
            bcd_2     : out std_logic_vector(6 downto 0)
        );
    end component;

begin
    -- Clock generation
    clk <= not clk after CLK_PERIOD/2 when not test_complete else '0';
    reset_n <= not reset;

    -- Unit Under Test
    uut: top
        port map (
            clk => clk,
            reset_n => reset_n,
            execute => execute,
            ms => ms,
            mr => mr,
            switch => switch,
            op => op,
            led => led,
            bcd_0 => bcd_0,
            bcd_1 => bcd_1,
            bcd_2 => bcd_2
        );

    -- Test process
    test_sequence: process
        procedure pulse_signal(signal sig: out std_logic; duration: in natural) is
        begin
            sig <= '1';
            for i in 1 to duration loop
                wait until rising_edge(clk);
            end loop;
            sig <= '0';
            wait until rising_edge(clk);
        end procedure;
        
        procedure wait_cycles(cycles: in natural) is
        begin
            for i in 1 to cycles loop
                wait until rising_edge(clk);
            end loop;
        end procedure;
        
        procedure check_result(expected: in integer; operation: in string) is
        begin
            wait_cycles(2); -- Allow result to propagate
            report "Operation: " & operation & " | Expected: " & integer'image(expected);
            -- Note: In simulation, we'd need to add signals to monitor internal results
        end procedure;

    begin
        -- Initialize
        report "Starting Calculator Test Bench";
        reset <= '1';
        wait_cycles(5);
        reset <= '0';
        wait_cycles(5);
        
        -- Test Sequence 1: Multiply 4 by 8
        report "Test 1: Multiply 4 by 8";
        switch <= std_logic_vector(to_unsigned(4, 8)); -- First operand (will be in working reg after reset)
        op <= "10"; -- Multiply operation
        wait_cycles(2);
        
        -- Load first operand (4) into working register (simulate initial state)
        -- Note: After reset, working register should be 0, so we need to set it
        switch <= std_logic_vector(to_unsigned(4, 8));
        pulse_signal(execute, 2);
        wait_cycles(5);
        
        -- Now multiply by 8
        switch <= std_logic_vector(to_unsigned(8, 8)); -- Second operand
        op <= "10"; -- Multiply
        pulse_signal(execute, 2);
        wait_cycles(10);
        check_result(32, "4 * 8 = 32");
        
        -- Test Sequence 2: Save result to memory
        report "Test 2: Save result (32) to memory";
        pulse_signal(ms, 2);
        wait_cycles(5);
        
        -- Test Sequence 3: Subtract 8
        report "Test 3: Subtract 8 from current value";
        switch <= std_logic_vector(to_unsigned(8, 8));
        op <= "01"; -- Subtract
        pulse_signal(execute, 2);
        wait_cycles(10);
        check_result(24, "32 - 8 = 24");
        
        -- Test Sequence 4: Divide by 2
        report "Test 4: Divide 24 by 2";
        switch <= std_logic_vector(to_unsigned(2, 8));
        op <= "11"; -- Divide
        pulse_signal(execute, 2);
        wait_cycles(10);
        check_result(12, "24 / 2 = 12");
        
        -- Test Sequence 5: Load saved number from memory
        report "Test 5: Load saved number (32) from memory";
        pulse_signal(mr, 2);
        wait_cycles(10);
        check_result(32, "Memory recall should give 32");
        
        -- Test Sequence 6: Divide saved number by 2
        report "Test 6: Divide saved number (32) by 2";
        switch <= std_logic_vector(to_unsigned(2, 8));
        op <= "11"; -- Divide
        pulse_signal(execute, 2);
        wait_cycles(10);
        check_result(16, "32 / 2 = 16");
        
        -- Final wait and completion
        wait_cycles(20);
        report "All test sequences completed successfully!";
        test_complete <= true;
        wait;
    end process;

    -- Monitor process to display internal state
    monitor: process
    begin
        wait until rising_edge(clk);
        if reset = '0' then
            report "Time: " & time'image(now) & 
                   " | LEDs: " & integer'image(to_integer(unsigned(led))) &
                   " | Op: " & integer'image(to_integer(unsigned(op))) &
                   " | Switches: " & integer'image(to_integer(unsigned(switch)));
        end if;
    end process;

end testbench;